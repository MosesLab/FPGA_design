-------------------------------------------------------------------------------
--$Date: 2007/08/01 23:10:49 $
--$RCSfile: example_tb_vhd.ejava,v $
--$Revision: 1.1.2.1 $
--------------------------------------------------------------------------------
--   ____  ____ 
--  /   /\/   / 
-- /___/  \  /    Vendor: Xilinx 
-- \   \   \/     Version : 1.7
--  \   \         Application : GTP Wizard 
--  /   /         Filename : example_tb.vhd
-- /___/   /\     Timestamp : 
-- \   \  /  \ 
--  \___\/\___\ 
--
--
-- Module EXAMPLE_TB
-- Generated by Xilinx GTP Wizard
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;
use work.ctiUtil.all;
use work.ctiSim.all;
use work.txt_util.all;

library modelsim_lib;
use modelsim_lib.util.all;

entity EXAMPLE_TB is
end EXAMPLE_TB;

architecture RTL of EXAMPLE_TB is

--*************************Parameter Declarations******************************

    constant   REFCLK_PERIOD        :   time :=  10.0 ns;
  
--**************************** Component Declarations *************************

    component mgt_tester 
    generic
    (
        EXAMPLE_SIM_GTPRESET_SPEEDUP    : integer    := 1;
        EXAMPLE_SIM_PLL_PERDIV2         : bit_vector := x"190";
        --EXAMPLE_USE_CHIPSCOPE           : integer    := 1     -- Set to 1 to use Chipscope to drive resets
			c_numgtp								: integer := 4
    );
    port
    (
    TILE0_REFCLK_PAD_N_IN                   : in   std_logic;
    TILE0_REFCLK_PAD_P_IN                   : in   std_logic;
	
    RXN_IN                                  : in   std_logic_vector(3 downto 0);
    RXP_IN                                  : in   std_logic_vector(3 downto 0);
    TXN_OUT                                 : out  std_logic_vector(3 downto 0);
    TXP_OUT                                 : out  std_logic_vector(3 downto 0);
	
	gtp_rst									: in std_logic;
	rx_rst 									: in std_logic;
	tx_rst 									: in std_logic;

	lb_clk									: in std_logic;
	lb_we									: in std_logic_vector(3 downto 0);
	lb_en									: in std_logic;
	lb_a									: in std_logic_vector(8 downto 2);
	lb_di									: in std_logic_vector(31 downto 0);
	lb_do									: out std_logic_vector(31 downto 0);
		
	lb_tx_start								: in std_logic_vector(3 downto 0);
	lb_tx_done								: out std_logic_vector(3 downto 0);
	lb_tx_sz								: in std_logic_vector(31 downto 0);
	
	lb_rx_done								: out std_logic_vector(3 downto 0);
	lb_rx_sz								: out std_logic_vector(31 downto 0);
	lb_rx_ok								: in std_logic_vector(3 downto 0);
	lb_rx_err_cnt							: out std_logic_vector(31 downto 0);
	
	lb_loopback								: in  std_logic_matrix_03(3 downto 0);
	tile0_pll_ok							: out std_logic;
	tile1_pll_ok							: out std_logic
	);
    end component mgt_tester;

    component SIM_RESET_MGT_MODEL 
    port 
    (
        GSR_IN     : in std_logic
    );
    end component;

--************************Internal Register Declarations***********************

--************************** Register Declarations ****************************        

    signal  debounce_pma_reset_r    :   std_logic_vector(0 to 3);
    signal  refclk_n_r              :   std_logic;
    signal  drp_clk_r               :   std_logic;
    signal  tx_usrclk_r             :   std_logic;
    signal  rx_usrclk_r             :   std_logic;    
    signal  gsr_r                   :   std_logic;
    signal  gts_r                   :   std_logic;
    signal  reset_i                 :   std_logic;

--********************************Wire Declarations**********************************
    
    ----------------------------------- Global Signals ------------------------------
    signal  refclk_p_r              :   std_logic;
    signal  tied_to_ground_i        :   std_logic;
    ---------------------------- Example Module Connections -------------------------
    signal  rxn_in_i                :   std_logic_vector(3 downto 0);
    signal  rxp_in_i                :   std_logic_vector(3 downto 0);
    signal  txn_out_i               :   std_logic_vector(3 downto 0);
    signal  txp_out_i               :   std_logic_vector(3 downto 0);

    signal  tile0_plllkdet_i       :   std_logic;
    signal  tile1_plllkdet_i       :   std_logic;

	-- MF signals
	signal connect : std_logic;

	signal t0ch0_framecheck_cnt : std_logic_vector(8 downto 0);
	signal t0ch0_framecheck_startchar : std_logic;	
	signal t0ch0_loopback : std_logic_vector(2 downto 0);
	signal simFinished : boolean  := false;
	
	
	--signal gtp_rst								:  std_logic;
	--signal rx_rst 								:  std_logic;
	--signal tx_rst 								:  std_logic;

	signal lb_clk								:  std_logic;
	signal lb_we								:  std_logic_vector(3 downto 0);
	signal lb_a									:  std_logic_vector(8 downto 2);
	signal lb_di								:  std_logic_vector(31 downto 0);
	signal lb_do								:  std_logic_vector(31 downto 0);
		
	signal lb_tx_start							:  std_logic_vector(3 downto 0);
	signal lb_tx_done							:  std_logic_vector(3 downto 0);
	signal lb_tx_sz								:  std_logic_vector(31 downto 0);
	
	signal lb_rx_done							:  std_logic_vector(3 downto 0);
	signal lb_rx_sz								:  std_logic_vector(31 downto 0);
	signal lb_rx_ok								:  std_logic_vector(3 downto 0);
	signal lb_rx_err_cnt						:  std_logic_vector(31 downto 0);
	
	signal lb_loopback							:  std_logic_matrix_03(3 downto 0); -- := (others => '0');
	signal tile0_pll_ok							:  std_logic;
	signal tile1_pll_ok							:  std_logic;	
	
	--signal pattern0 :      std_logic_matrix_08(0 to 127);

	constant c_sz_buf : integer := 16;  -- 16 *32 = 512 bits
	
	
--*********************************Main Body of Code**********************************
begin

    -- ------------------------------- Tie offs -------------------------------   
    tied_to_ground_i        <=  '0';
    
    -- ------------------------- MGT Serial Connections -----------------------
    rxn_in_i                <=  txn_out_i when connect='1' else (others=>'0');
    rxp_in_i                <=  txp_out_i when connect='1' else (others=>'1');  

    ------- Instantiate the ROC module for resetting the VHDL MGT Smart Model ------
    sim_reset_mgt_model_i : SIM_RESET_MGT_MODEL  
    port map    
    (
        GSR_IN           =>           reset_i
    );

    ---------------------- Generate Reference Clock input  --------------------
    process
    begin
        refclk_n_r  <=  '1';
        wait for REFCLK_PERIOD/2;
        refclk_n_r  <=  '0';
        wait for REFCLK_PERIOD/2;
    end process;

    refclk_p_r <= not refclk_n_r;
	
	process
	begin
		lb_clk <= '1';
		wait for 10 ns;
		lb_clk <= '0';
		wait for 10 ns;
	end process;
                      
    ----------------------------------- Resets ---------------------------------
    --process
    --begin
    --    reset_i <= '1';
    --    wait for 100 ns;
     --   reset_i <= '0';
     --   wait; 
    --end process;

    ------------------- Instantiate an EXAMPLE_MGT_TOP module  -----------------
    example_mgt_top_i : mgt_tester
    generic map
    (
        EXAMPLE_SIM_GTPRESET_SPEEDUP        =>  1,        -- Speedup is turned on for simulation
        EXAMPLE_SIM_PLL_PERDIV2             =>  x"1f4"      -- Set to the VCO Unit Interval time
											-- was x190

    )
    port map
    (
        TILE0_REFCLK_PAD_N_IN       =>  refclk_n_r,   
        TILE0_REFCLK_PAD_P_IN       =>  refclk_p_r,

        RXN_IN                      =>  rxn_in_i,
        RXP_IN                      =>  rxp_in_i,
        TXN_OUT                     =>  txn_out_i,
        TXP_OUT                     =>  txp_out_i,

		gtp_rst						=> reset_i,
		rx_rst 						=> '0',
		tx_rst 						=> '0',

		lb_clk						=> lb_clk,
		lb_we						=> lb_we,
		lb_en						=> '1',
		lb_a						=> lb_a,
		lb_di						=> lb_di,
		lb_do						=> lb_do,
			
		lb_tx_start					=> lb_tx_start,
		lb_tx_done					=> lb_tx_done,
		lb_tx_sz					=> lb_tx_sz,
		
		lb_rx_done					=> lb_rx_done,
		lb_rx_sz					=> lb_rx_sz,
		lb_rx_ok					=> lb_rx_ok,
		lb_rx_err_cnt				=> lb_rx_err_cnt,
		
		lb_loopback					=> lb_loopback,
		tile0_pll_ok				=> tile0_plllkdet_i,
		tile1_pll_ok				=> tile1_plllkdet_i
    );

    ------------------------------------
	
	-- signal spy
	
    -- spy_process : process
	-- begin
        -- init_signal_spy("/example_tb/example_mgt_top_i/tile0_frame_check0/rx_data_has_start_char_c","/EXAMPLE_TB/t0ch0_framecheck_startchar",1,1);	
        -- init_signal_spy("/example_tb/example_mgt_top_i/tile0_frame_check0/read_counter_i","/EXAMPLE_TB/t0ch0_framecheck_cnt",1,1);
        -- wait;
    -- end process spy_process;
	
	-- spy_enable_disable : process
	-- begin
		-- wait for 1 ns;
        -- enable_signal_spy("/example_tb/example_mgt_top_i/tile0_frame_check0/rx_data_has_start_char_c","/EXAMPLE_TB/t0ch0_framecheck_startchar",0);			
        -- enable_signal_spy("/example_tb/example_mgt_top_i/tile0_frame_check0/read_counter_i","/EXAMPLE_TB/t0ch0_framecheck_cnt",0);
		-- wait;
    -- end process spy_enable_disable;
        
	--drive_sig_process : process
	--begin
	--	init_signal_driver("/EXAMPLE_TB/t0ch0_loopback", "/example_tb/example_mgt_top_i/pciegtp_wrapper_i/tile0_pciegtp_wrapper_i/loopback0_in", open, open, 1);
	--	wait;
	--end process drive_sig_process;	
	
	tests : process
	
		procedure writeBuffer(num : integer; tx_or_rx : std_logic; pat : std_logic_matrix_32) is
		begin
		
			wait until rising_edge(lb_clk);
			wait for 3 ns;
			lb_di <= x"00000000";
			lb_we <= x"0";
				
			for i in 0 to (c_sz_buf-1) loop	
				wait until rising_edge(lb_clk);
				wait for 3 ns;
				lb_a(8) <= tx_or_rx;
				lb_a(7 downto 6) <= std_logic_vector( to_unsigned(num,2) );
				lb_a(5 downto 2) <= std_logic_vector( to_unsigned(i,4) );
				lb_we <= x"F";
				lb_di <= pat(i);
			end loop;

			wait until rising_edge(lb_clk);
			wait for 3 ns;
			lb_di <= x"00000000";
			lb_we <= x"0";
		end procedure;
		
		procedure verifyBuffer(num : integer; tx_or_rx : std_logic; pat : std_logic_matrix_32) is
		begin
			wait until rising_edge(lb_clk);		
			
			for i in 0 to (c_sz_buf-1) loop
				wait for 1 ns;
				lb_a(8) <= tx_or_rx;
				lb_a(7 downto 6) <= std_logic_vector( to_unsigned(num,2) );
				lb_a(5 downto 2) <= std_logic_vector( to_unsigned(i,4) );
				
				wait until rising_edge(lb_clk);
				wait for 3 ns;
				assert (lb_do  = pat(i))
	            	report "buffer does not match @ " & str(i) & " Expected " & hstr(pat(i)) & " Read " & hstr(lb_do)
				    severity failure;		   
			end loop;
		end procedure;

		variable pat_clr : std_logic_matrix_32(0 to (c_sz_buf-1));
		variable pat_0 : std_logic_matrix_32(0 to (c_sz_buf-1));
		variable done_mask : std_logic_vector(3 downto 0);
	begin
	   title("Simulation starting");
	   lb_loopback(0) <= "000";
	   lb_loopback(1) <= "000";
	   lb_loopback(2) <= "000";
	   lb_loopback(3) <= "000";
	   
		lb_we  <= (others => '0');
		lb_a  <= (others => '0');
		lb_tx_start  <= (others => '0');
		lb_tx_sz  <= (others => '0');
		lb_rx_sz  <= (others => '0');
		lb_rx_ok <= (others => '0');	  

		for i in 0 to (c_sz_buf-1) loop
			pat_clr(i) := (others => '0');
		end loop;
		
	    connect <= '1';
	    --t0ch0_loopback <= "000";

		wait for 10 ns;
		
		reset_i <= '1';
        wait for 100 ns;
        reset_i <= '0';
		
		msg("Reset done");
		
		
		
		while tile0_plllkdet_i /= '1' loop
			wait for 100 ns;	
			msg("Waiting for PLL ready");
		end loop;
		
		msg("PLL ready");
	
	for gtp in 0 to 3 loop
		title("testing gtp #" & str(gtp));
	
		msg("clearing tx buffer" );
		writeBuffer(gtp,'0',pat_clr);
		
		msg("clearing rx buffer");
		writeBuffer(gtp,'1',pat_clr);
		
		msg("verify tx buffer empty");
		verifyBuffer(gtp, '0', pat_clr);
		
		msg("verify rx buffer empty");
		verifyBuffer(gtp, '1', pat_clr);
		
		wait for 100 ns;

		msg("Generate pat_0");
		
		for i in 0 to (c_sz_buf-1) loop
			pat_0(i)(7 downto 0) := std_logic_vector( to_unsigned(i*4+0,8) );
			pat_0(i)(1 downto 0) := std_logic_vector( to_unsigned(gtp,2) );
			pat_0(i)(15 downto 8) := std_logic_vector( to_unsigned(i*4+1,8) );
			pat_0(i)(23 downto 16) := std_logic_vector( to_unsigned(i*4+2,8) );
			pat_0(i)(31 downto 24) := std_logic_vector( to_unsigned(i*4+3,8) );
		end loop;	

		pat_0(0)(7 downto 0) := x"FF";
		

		msg("writing to tx buffer");
		writeBuffer(gtp,'0',pat_0);
			
		msg("verifying tx buffer");
		verifyBuffer(gtp, '0', pat_0);		
		
		wait until rising_edge(lb_clk);
		wait for 2 ns;
		msg("Enable receiver");
		lb_rx_ok(gtp) <= '1';
		lb_tx_sz <= x"00000000";
		lb_tx_sz(7+gtp*8 downto gtp*8) <= x"3F"; --64 (size in bytes)
		
		wait until rising_edge(lb_clk);
		wait for 2 ns;
		msg("start transmitter");
		lb_tx_start(gtp) <= '1';
		
		done_mask := "0000";
		done_mask(gtp) := '1';
		
		while (lb_tx_done /= done_mask) loop
			wait for 50 ns;	
			msg("Waiting for tx done");
		end loop;
		
		lb_tx_start(gtp) <= '0';		
		
		while lb_rx_done /= done_mask loop
			wait for 50 ns;	
			msg("Waiting for rx done");
		end loop;
				
		msg("clearing tx buffer ");
		writeBuffer(gtp,'0',pat_clr);
		
		msg("verify rx buffer has pat_0");
		verifyBuffer(gtp, '1', pat_0);		
		

		lb_rx_ok(gtp) <= '0';
	
		wait for 500 ns;
	end loop;
	
		-- wait until t0ch0_framecheck_startchar = '1';
		-- msg("Hit start character");
		
		-- wait until t0ch0_framecheck_cnt = to_stdlogic(16#10#,9);

		-- msg("Frame check hit 0x10");
		-- msg("Disconnecting");		
		-- connect <= '0';
		-- wait for 100 ns;

		-- msg("Reconnecting");				
		-- connect <= '1';		

		-- wait for 1 us;
		
		
		-- msg("Change loopback mode - near end PCS (001)");
		-- connect <= '0';
		-- t0ch0_loopback <= "001";
		
        -- reset_i <= '1';
        -- wait for 100 ns;
        -- reset_i <= '0';

		-- wait for 100 ns;	
		-- wait until tile0_plllkdet_i = '1';
		-- msg("PLL ready");
		
		--signal_force("/example_tb/example_mgt_top_i/pciegtp_wrapper_i/tile0_pciegtp_wrapper_i/loopback0_in", "001", 0 ns, drive, open, 1);		
		-- wait for 1 us;
		
		-- msg("Change loopback mode - near end PMA (010)");
		-- t0ch0_loopback <= "010";
		
        -- reset_i <= '1';
        -- wait for 100 ns;
        -- reset_i <= '0';
		
		-- wait for 100 ns;	
		-- wait until tile0_plllkdet_i = '1';
		-- msg("PLL ready");		
		
		--signal_force("/example_tb/example_mgt_top_i/pciegtp_wrapper_i/tile0_pciegtp_wrapper_i/loopback0_in", "010", 0 ns, drive, open, 1);				
		-- wait for 1 us;
		
		title("Finished");
		simFinished <= TRUE;
		
		wait;
	
	end process;
	
end RTL;

